module main

// TODO
