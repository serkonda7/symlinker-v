module linker
